module Hello2(
);
	initial begin
		$display("Hello,World");
	end
endmodule	
