module Hello (
	);
	initial begin
		$display("Hello,World");
		$display("wktk");
	end
endmodule
